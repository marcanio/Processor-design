library IEEE;
use IEEE.std_logic_1164.all;

entity Decoder5to32 is
 generic(N : integer := 32);
  port(input5           : in std_logic_vector(4 downto 0);     -- 5 Bit input
       output32         : out std_logic_vector(31 downto 0);
       enable		: in std_logic);   -- Enable bit

end Decoder5to32;


architecture DataFlow of Decoder5to32 is

begin

process(input5, enable)
begin
	output32 <= "00000000000000000000000000000000"; --Default output
	
	if (enable = '1') then
		case input5 is
			when "00000" => output32 <= "00000000000000000000000000000001";
			when "00001" => output32 <= "00000000000000000000000000000010";
			when "00010" => output32 <= "00000000000000000000000000000100";	
			when "00011" => output32 <= "00000000000000000000000000001000";	
			when "00100" => output32 <= "00000000000000000000000000010000";
			when "00101" => output32 <= "00000000000000000000000000100000";
			when "00110" => output32 <= "00000000000000000000000001000000";
			when "00111" => output32 <= "00000000000000000000000010000000";
			when "01000" => output32 <= "00000000000000000000000100000000";	
			when "01001" => output32 <= "00000000000000000000001000000000";	
			when "01010" => output32 <= "00000000000000000000010000000000"; 
			when "01011" => output32 <= "00000000000000000000100000000000";
			when "01100" => output32 <= "00000000000000000001000000000000";
			when "01101" => output32 <= "00000000000000000010000000000000";
			when "01110" => output32 <= "00000000000000000100000000000000";	
			when "01111" => output32 <= "00000000000000001000000000000000";	
			when "10000" => output32 <= "00000000000000010000000000000000";
			when "10001" => output32 <= "00000000000000100000000000000000";
			when "10010" => output32 <= "00000000000001000000000000000000";
			when "10011" => output32 <= "00000000000010000000000000000000";
			when "10100" => output32 <= "00000000000100000000000000000000";	
			when "10101" => output32 <= "00000000001000000000000000000000";	
			when "10110" => output32 <= "00000000010000000000000000000000";
			when "10111" => output32 <= "00000000100000000000000000000000";
			when "11000" => output32 <= "00000001000000000000000000000000";
			when "11001" => output32 <= "00000010000000000000000000000000";
			when "11010" => output32 <= "00000100000000000000000000000000";	
			when "11011" => output32 <= "00001000000000000000000000000000";	
			when "11100" => output32 <= "00010000000000000000000000000000";
			when "11101" => output32 <= "00100000000000000000000000000000";
			when "11110" => output32 <= "01000000000000000000000000000000";
			when "11111" => output32 <= "10000000000000000000000000000000";
			when others  => output32 <= "00000000000000000000000000000000";
		end case;
	end if;
end process;
end DataFlow;









